module WallaceTree (
		                   input  wire [11:0] A,
                       input  wire [11:0] B,
		                   output wire [23:0] M
                   );

  wire S[135:0];
  wire C[139:0];

  // M[ 0] : 1
  assign M[0] = B[0] & A[0];

  // M[ 1] : 2
  FA m0 ( B[ 0]&A[ 1] , B[ 1]&A[ 0] ,        1'b0 , M[ 1] , C[ 0] );

  // M[ 2] : 3
  FA m1 ( B[ 0]&A[ 2] , B[ 1]&A[ 1] , B[ 2]&A[ 0] , S[ 0] , C[ 1] );

  FA m2 (       S[ 0] ,       C[ 0] ,        1'b0 , M[ 2] , C[ 2] );

  // M[ 3] : 4
  FA m3 ( B[ 0]&A[ 3] , B[ 1]&A[ 2] , B[ 2]&A[ 1] , S[ 1] , C[ 3] );

  FA m4 (       S[ 1] ,       C[ 1] , B[ 3]&A[ 0] , S[ 2] , C[ 4] );

  FA m5 (       S[ 2] ,       C[ 2] ,        1'b0 , M[ 3] , C[ 5] );                       

  // M[ 4] : 5
  FA m6 ( B[ 0]&A[ 4] , B[ 1]&A[ 3] , B[ 2]&A[ 2] , S[ 3] , C[ 6] );
  FA m7 (        1'b0 , B[ 3]&A[ 1] , B[ 4]&A[ 0] , S[ 4] , C[ 7] );

  FA m8 (       S[ 3] ,       S[ 4] ,       C[ 3] , S[ 5] , C[ 8] );

  FA m9 (       S[ 5] ,        1'b0 ,       C[ 4] , S[ 6] , C[ 9] ); 

  FA m10(       S[ 6] ,        1'b0 ,       C[ 5] , M[ 4] , C[10] );       

  // M[ 5] : 6
  FA m11( B[ 0]&A[ 5] , B[ 1]&A[ 4] , B[ 2]&A[ 3] , S[ 7] , C[11] );
  FA m12( B[ 3]&A[ 2] , B[ 4]&A[ 1] , B[ 5]&A[ 0] , S[ 8] , C[12] );

  FA m13(       S[ 7] ,       C[ 6] ,       C[ 7] , S[ 9] , C[13] );

  FA m14(       S[ 8] ,       S[ 9] ,       C[ 8] , S[10] , C[14] );

  FA m15(       S[10] ,        1'b0 ,       C[ 9] , S[11] , C[15] ); 

  FA m16(       S[11] ,        1'b0 ,       C[10] , S[12] , C[16] );

  // M[ 6] : 7
  FA m17( B[ 0]&A[ 6] , B[ 1]&A[ 5] , B[ 2]&A[ 4] , S[13] , C[17] );
  FA m18( B[ 3]&A[ 3] , B[ 4]&A[ 2] , B[ 5]&A[ 1] , S[14] , C[18] );

  FA m19(       S[13] ,       S[14] , B[ 6]&A[ 0] , S[15] , C[19] );
  FA m20(       C[11] ,       C[12] ,        1'b0 , S[16] , C[20] );
  
  FA m21(       S[15] ,       S[16] ,       C[14] , S[17] , C[21] );

  FA m22(       S[17] ,       C[15] ,        1'b0 , S[18] , C[22] ); 

  FA m23(       S[18] ,       C[16] ,        1'b0 , S[19] , C[23] );

  // M[ 7] : 8

  FA m24( B[ 0]&A[ 7] , B[ 1]&A[ 6] , B[ 2]&A[ 5] , S[20] , C[24] );
  FA m25( B[ 3]&A[ 4] , B[ 4]&A[ 3] , B[ 5]&A[ 2] , S[21] , C[25] );
  FA m26( B[ 6]&A[ 1] , B[ 7]&A[ 0] ,        1'b0 , S[22] , C[26] );

  FA m27(       S[20] ,       S[21] ,       S[22] , S[23] , C[27] );
  FA m28(       C[17] ,       C[18] ,        1'b0 , S[24] , C[28] );

  FA m29(       S[23] ,       S[24] ,       C[19] , S[25] , C[29] );
  
  FA m30(       S[25] ,       C[20] ,       C[21] , S[26] , C[30] );
 
  FA m31(       S[26] ,       C[22] ,        1'b0 , S[27] , C[31] );

 
  // M[ 8] : 9            
  FA m32( B[ 0]&A[ 8] , B[ 1]&A[ 7] , B[ 2]&A[ 6] , S[28] , C[32] );
  FA m33( B[ 3]&A[ 5] , B[ 4]&A[ 4] , B[ 5]&A[ 3] , S[29] , C[33] );
  FA m34( B[ 6]&A[ 2] , B[ 7]&A[ 1] , B[ 8]&A[ 0] , S[30] , C[34] );

  FA m35(       S[28] ,       S[29] ,       S[30] , S[31] , C[35] );
  FA m36(       C[24] ,       C[25] ,       C[26] , S[32] , C[36] );

  FA m37(       S[31] ,       S[32] ,       C[27] , S[33] , C[37] );

  FA m38(       S[33] ,       C[28] ,       C[29] , S[34] , C[38] );
  
  FA m39(       S[34] ,       C[30] ,        1'b0 , S[35] , C[39] );

  
  // M[ 9] : 10
  FA m40( B[ 0]&A[ 9] , B[ 1]&A[ 8] , B[ 2]&A[ 7] , S[36] , C[40] );
  FA m41( B[ 3]&A[ 6] , B[ 4]&A[ 5] , B[ 5]&A[ 4] , S[37] , C[41] );
  FA m42( B[ 6]&A[ 3] , B[ 7]&A[ 2] , B[ 8]&A[ 1] , S[38] , C[42] );

  FA m43(       S[36] ,       S[37] ,       S[38] , S[39] , C[43] );
  FA m44(       C[32] ,       C[33] ,       C[34] , S[40] , C[44] );

  FA m45(       S[39] ,       S[40] , B[ 9]&A[ 0] , S[41] , C[45] );
  FA m46(       C[35] ,       C[36] ,        1'b0 , S[42] , C[46] );
  
  FA m47(       S[41] ,       S[42] ,       C[37] , S[43] , C[47] );

  FA m48(       S[43] ,       C[38] ,        1'b0 , S[44] , C[48] );

           
  // M[10] : 11
  FA m49( B[ 0]&A[10] , B[ 1]&A[ 9] , B[ 2]&A[ 8] , S[45] , C[49] );
  FA m50( B[ 3]&A[ 7] , B[ 4]&A[ 6] , B[ 5]&A[ 5] , S[46] , C[50] ); 
  FA m51( B[ 6]&A[ 4] , B[ 7]&A[ 3] , B[ 8]&A[ 2] , S[47] , C[51] );
  FA m52( B[ 9]&A[ 1] , B[10]&A[ 0] ,        1'b0 , S[48] , C[52] );

  FA m53(       S[44] ,       S[45] ,       S[46] , S[49] , C[53] );
  FA m54(       C[40] ,       C[41] ,       C[42] , S[50] , C[54] );

  FA m55(       S[48] ,       S[49] ,       S[50] , S[51] , C[55] );
  FA m56(       C[43] ,       C[44] ,        1'b0 , S[52] , C[56] );

  FA m57(       S[51] ,       S[52] ,       C[45] , S[53] , C[57] ); 

  FA m58(       S[53] ,       C[46] ,       C[47] , S[54] , C[58] ); 

  
  // M[11] : 12
  FA m59( B[ 0]&A[11] , B[ 1]&A[10] , B[ 2]&A[ 9] , S[55] , C[59] );
  FA m60( B[ 3]&A[ 8] , B[ 4]&A[ 7] , B[ 5]&A[ 6] , S[56] , C[60] );
  FA m61( B[ 6]&A[ 5] , B[ 7]&A[ 4] , B[ 8]&A[ 3] , S[57] , C[61] );
  FA m62( B[ 9]&A[ 2] , B[10]&A[ 1] , B[11]&A[ 0] , S[58] , C[62] );

  FA m63(       C[49] ,       C[50] ,       C[51] , S[59] , C[63] );
  FA m64(       S[55] ,       S[56] ,       S[57] , S[60] , C[64] );
  FA m65(       C[52] ,       S[58] ,        1'b0 , S[61] , C[65] );
  
  FA m66(       S[59] ,       S[60] ,       S[61] , S[62] , C[66] );
  FA m67(       C[53] ,       C[54] ,        1'b0 , S[63] , C[67] );

  FA m68(       S[62] ,       S[63] ,       C[55] , S[64] , C[68] );

  FA m69(       S[64] ,       C[56] ,       C[57] , S[65] , C[69] );

  
  // M[12] : 11
  FA m70( B[ 1]&A[11] , B[ 2]&A[10] ,        1'b0 , S[66] , C[70] );
  FA m71( B[ 3]&A[ 9] , B[ 4]&A[ 8] , B[ 5]&A[ 7] , S[67] , C[71] );
  FA m72( B[ 6]&A[ 6] , B[ 7]&A[ 5] , B[ 8]&A[ 4] , S[68] , C[72] );
  FA m73( B[ 9]&A[ 3] , B[10]&A[ 2] , B[11]&A[ 1] , S[69] , C[73] );

  FA m74(       C[59] ,       C[60] ,       C[61] , S[70] , C[74] );
  FA m75(       S[66] ,       S[67] ,       S[68] , S[71] , C[75] );
  FA m76(       C[62] ,       S[69] ,        1'b0 , S[72] , C[76] );

  FA m77(       C[63] ,       C[64] ,       C[65] , S[73] , C[77] );
  FA m78(       C[70] ,       C[71] ,       C[72] , S[74] , C[78] ); 

  FA m79(       S[73] ,       S[74] ,       C[66] , S[75] , C[79] );

  FA m80(       S[75] ,       C[67] ,       C[68] , S[76] , C[80] );


  // M[13] : 10
  FA m81( B[ 3]&A[10] , B[ 4]&A[ 9] , B[ 5]&A[ 8] , S[77] , C[81] );
  FA m82( B[ 6]&A[ 7] , B[ 7]&A[ 6] , B[ 8]&A[ 5] , S[78] , C[82] );
  FA m83( B[ 9]&A[ 4] , B[10]&A[ 3] , B[11]&A[ 2] , S[79] , C[83] );

  FA m84(       S[77] ,       S[78] ,       S[79] , S[80] , C[84] );
  FA m85(       C[70] ,       C[71] ,       C[72] , S[81] , C[85] );
  FA m86(       C[73] , B[ 2]&A[11] ,        1'b0 , S[82] , C[86] );

  FA m87(       C[74] ,       C[75] ,       C[76] , S[83] , C[87] );
  FA m88(       S[80] ,       S[81] ,       S[82] , S[84] , C[88] );

  FA m89(       S[83] ,       S[84] ,       C[77] , S[85] , C[89] );

  FA m90(       S[85] ,       C[78] ,       C[79] , S[86] , C[90] );
  
                   
  // M[14] : 9
  FA m91( B[ 3]&A[11] , B[ 4]&A[10] , B[ 5]&A[ 9] , S[87] , C[91] );
  FA m92( B[ 6]&A[ 8] , B[ 7]&A[ 7] , B[ 8]&A[ 6] , S[88] , C[92] );
  FA m93( B[ 9]&A[ 5] , B[10]&A[ 4] , B[11]&A[ 3] , S[89] , C[93] );

  FA m94(       S[87] ,       S[88] ,       S[89] , S[90] , C[94] );
  FA m95(       C[81] ,       C[82] ,       C[83] , S[91] , C[95] );

  FA m96(       C[84] ,       C[85] ,       C[86] , S[92] , C[96] );
  FA m97(       S[90] ,       S[91] ,        1'b0 , S[93] , C[97] );

  FA m98(       S[92] ,       S[93] ,       C[87] , S[94] , C[98] );

  FA m99(       S[94] ,       C[88] ,       C[89] , S[95] , C[99] );

     
  // M[15] : 8
  FA m100(B[ 4]&A[11] , B[ 5]&A[10] ,        1'b0 , S[96] , C[100]);
  FA m101(B[ 6]&A[ 9] , B[ 7]&A[ 8] , B[ 8]&A[ 7] , S[97] , C[101]);
  FA m102(B[ 9]&A[ 6] , B[10]&A[ 5] , B[11]&A[ 4] , S[98] , C[102]);

  FA m103(      S[96] ,       S[97] ,       S[98] , S[99] , C[103]);
  FA m104(      C[91] ,       C[92] ,       C[93] , S[100], C[104]);

  FA m105(      S[99] ,       S[100],       C[94] , S[101], C[105]);

  FA m106(      S[101],       C[95] ,       C[96] , S[102], C[106]);

  FA m107(      S[102],       C[97] ,       C[98] , S[103], C[107]);

         
  // M[16] : 7
  FA m108(B[ 6]&A[10] , B[ 7]&A[ 9] , B[ 8]&A[ 8] , S[104], C[108]);
  FA m109(B[ 9]&A[ 7] , B[10]&A[ 6] , B[11]&A[ 5] , S[105], C[109]);

  FA m110(      S[104],      S[105] , B[ 5]&A[11] , S[106], C[110]);
  FA m111(      C[100],      C[101] ,      C[102] , S[107], C[111]);

  FA m112(      S[106],      S[107] ,      C[103] , S[108], C[112]);

  FA m113(      S[108],      C[104] ,      C[105] , S[109], C[113]);

  FA m114(      S[109],      C[106] ,        1'b0 , S[110], C[114]);

  
  // M[17] : 6
  FA m115(B[ 6]&A[11] , B[ 7]&A[10] , B[ 8]&A[ 9] , S[111], C[115]);
  FA m116(B[ 9]&A[ 8] , B[10]&A[ 7] , B[11]&A[ 6] , S[112], C[116]);
  
  FA m117(      S[111],      S[112],       C[108] , S[113], C[117]);

  FA m118(      S[113],      C[109],       C[110] , S[114], C[118]);

  FA m119(      S[114],      C[111],       C[112] , S[115], C[119]);
 
  FA m120(      S[115],      C[113],         1'b0 , S[116], C[120]);


  // M[18] : 5
  FA m121(B[ 7]&A[11] , B[ 8]&A[10] ,        1'b0 , S[117], C[121]);
  FA m122(B[ 9]&A[ 9] , B[10]&A[ 8] , B[11]&A[ 7] , S[118], C[122]); 

  FA m123(     S[117] ,      S[118] ,      C[115] , S[119], C[123]);
  
  FA m124(     S[119] ,      C[116] ,      C[117] , S[120], C[124]);

  FA m125(     S[120] ,      C[118] ,        1'b0 , S[121], C[125]);        
  
  FA m126(     S[121] ,      C[119] ,        1'b0 , S[122], C[126]);

 
  // M[19] : 4
  FA m127(B[ 9]&A[10] , B[10]&A[ 9] , B[11]&A[ 8] , S[123], C[127]);
  
  FA m128(B[ 8]&A[11] ,      S[123] ,      C[121] , S[124], C[128]);

  FA m129(     S[124] ,      C[122] ,      C[123] , S[125], C[129]);

  FA m130(     S[125] ,      C[124] ,        1'b0 , S[126], C[130]);

  FA m131(     S[126] ,      C[125] ,        1'b0 , S[127], C[131]);
    

  // M[20] : 3
  FA m132(B[ 9]&A[11] , B[10]&A[10] , B[11]&A[ 9] , S[128], C[132]);

  // Nothing in level 2

  FA m133(     S[128] ,      C[127] ,      C[128] , S[129], C[133]);

  FA m134(     S[129] ,      C[129] ,        1'b0 , S[130], C[134]);

  FA m135(     S[130] ,      C[130] ,        1'b0 , S[131], C[135]);


  // M[21] : 2
  // Nothing in level 1

  FA m136(B[10]&A[11] , B[11]&A[10] ,      C[132] , S[132], C[136]);

  // Nothing in level 3

  FA m137(     S[132] ,      C[133] ,        1'b0 , S[133], C[137]);

  FA m138(     S[133] ,      C[134] ,        1'b0 , S[134], C[138]);


  // M[22] : 1
  // Just level 5
  FA m139(     S[134] ,      C[136] ,      C[137] , S[135], C[139]);


  assign M[23:5] = {C[139],C[138],C[135],C[131],C[126],C[120],C[114],C[107],C[99],C[90],C[80],C[69],C[58],C[48],C[39],C[31],C[23],C[16],C[10]}
                + { 1'b0,S[135],S[134],S[131],S[127],S[122],S[116],S[110],S[103],S[95],S[86],S[76],S[65],S[54],S[44],S[35],S[27],S[19],C[12]}; 
    

endmodule


module FA(
            // Inputs
            input  wire A,
            input  wire B,
            input  wire Cin,
            // Outputs
            output wire S,
            output wire Cout
         );
 
 assign {Cout,S}=A+B+Cin;

endmodule
